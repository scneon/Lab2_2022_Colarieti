library verilog;
use verilog.vl_types.all;
entity ParteA_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ParteA_vlg_check_tst;
