-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 25 03:30:55 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ParteD IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z0 : OUT STD_LOGIC;
        Z1 : OUT STD_LOGIC;
        Z2 : OUT STD_LOGIC;
        Z3 : OUT STD_LOGIC
    );
END ParteD;

ARCHITECTURE BEHAVIOR OF ParteD IS
    TYPE type_fstate IS (I,A1,B1,A2,B2,A3,B3,B4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= I;
            Z0 <= '0';
            Z1 <= '0';
            Z2 <= '0';
            Z3 <= '0';
        ELSE
            Z0 <= '0';
            Z1 <= '0';
            Z2 <= '0';
            Z3 <= '0';
            CASE fstate IS
                WHEN I =>
                    IF ((x = '0')) THEN
                        reg_fstate <= A1;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= I;
                    END IF;

                    Z3 <= '0';

                    Z2 <= '0';

                    Z1 <= '0';

                    Z0 <= '0';
                WHEN A1 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= A2;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A1;
                    END IF;

                    Z3 <= '0';

                    Z2 <= '1';

                    Z1 <= '1';

                    Z0 <= '0';
                WHEN B1 =>
                    reg_fstate <= B2;

                    Z3 <= '1';

                    Z2 <= '0';

                    Z1 <= '0';

                    Z0 <= '0';
                WHEN A2 =>
                    reg_fstate <= A3;

                    Z3 <= '1';

                    Z2 <= '1';

                    Z1 <= '1';

                    Z0 <= '1';
                WHEN B2 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B3;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= A2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B2;
                    END IF;

                    Z3 <= '1';

                    Z2 <= '1';

                    Z1 <= '0';

                    Z0 <= '0';
                WHEN A3 =>
                    reg_fstate <= I;

                    Z3 <= '1';

                    Z2 <= '0';

                    Z1 <= '1';

                    Z0 <= '1';
                WHEN B3 =>
                    reg_fstate <= B4;

                    Z3 <= '1';

                    Z2 <= '1';

                    Z1 <= '1';

                    Z0 <= '1';
                WHEN B4 =>
                    reg_fstate <= I;

                    Z3 <= '1';

                    Z2 <= '1';

                    Z1 <= '0';

                    Z0 <= '0';
                WHEN OTHERS => 
                    Z0 <= 'X';
                    Z1 <= 'X';
                    Z2 <= 'X';
                    Z3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
