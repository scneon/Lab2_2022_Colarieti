-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Nov 25 02:51:24 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Block1 IS 
	PORT
	(
		CLOCK :  IN  STD_LOGIC;
		SR :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		S0 :  OUT  STD_LOGIC;
		S1 :  OUT  STD_LOGIC;
		S2 :  OUT  STD_LOGIC;
		S3 :  OUT  STD_LOGIC;
		S :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC;
		V :  OUT  STD_LOGIC;
		C :  OUT  STD_LOGIC
	);
END Block1;

ARCHITECTURE bdf_type OF Block1 IS 

COMPONENT parteb_ffd
	PORT(D : IN STD_LOGIC;
		 CLOCK : IN STD_LOGIC;
		 Q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sumador_completo
	PORT(a : IN STD_LOGIC;
		 b : IN STD_LOGIC;
		 cin : IN STD_LOGIC;
		 f : OUT STD_LOGIC;
		 cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;


BEGIN 
S0 <= SYNTHESIZED_WIRE_31;
S1 <= SYNTHESIZED_WIRE_33;
S2 <= SYNTHESIZED_WIRE_32;
S3 <= SYNTHESIZED_WIRE_36;
S <= SYNTHESIZED_WIRE_36;



SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1 AND SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38;


b2v_DA0 : parteb_ffd
PORT MAP(D => A0,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_10);


b2v_DA1 : parteb_ffd
PORT MAP(D => A1,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_12);


b2v_DA2 : parteb_ffd
PORT MAP(D => A2,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_15);


b2v_DA3 : parteb_ffd
PORT MAP(D => A3,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_37);


b2v_DB0 : parteb_ffd
PORT MAP(D => B0,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_27);


b2v_DB1 : parteb_ffd
PORT MAP(D => B1,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_28);


b2v_DB2 : parteb_ffd
PORT MAP(D => B2,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_29);


b2v_DB3 : parteb_ffd
PORT MAP(D => B3,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_38);


b2v_DS0 : parteb_ffd
PORT MAP(D => SYNTHESIZED_WIRE_6,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_31);


b2v_DS1 : parteb_ffd
PORT MAP(D => SYNTHESIZED_WIRE_7,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_33);


b2v_DS2 : parteb_ffd
PORT MAP(D => SYNTHESIZED_WIRE_8,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_32);


b2v_DS3 : parteb_ffd
PORT MAP(D => SYNTHESIZED_WIRE_9,
		 CLOCK => CLOCK,
		 Q => SYNTHESIZED_WIRE_36);


b2v_FA0 : sumador_completo
PORT MAP(a => SYNTHESIZED_WIRE_10,
		 b => SYNTHESIZED_WIRE_11,
		 cin => SR,
		 f => SYNTHESIZED_WIRE_6,
		 cout => SYNTHESIZED_WIRE_14);


b2v_FA1 : sumador_completo
PORT MAP(a => SYNTHESIZED_WIRE_12,
		 b => SYNTHESIZED_WIRE_13,
		 cin => SYNTHESIZED_WIRE_14,
		 f => SYNTHESIZED_WIRE_7,
		 cout => SYNTHESIZED_WIRE_17);


b2v_FA2 : sumador_completo
PORT MAP(a => SYNTHESIZED_WIRE_15,
		 b => SYNTHESIZED_WIRE_16,
		 cin => SYNTHESIZED_WIRE_17,
		 f => SYNTHESIZED_WIRE_8,
		 cout => SYNTHESIZED_WIRE_20);


b2v_FA3 : sumador_completo
PORT MAP(a => SYNTHESIZED_WIRE_37,
		 b => SYNTHESIZED_WIRE_19,
		 cin => SYNTHESIZED_WIRE_20,
		 f => SYNTHESIZED_WIRE_9,
		 cout => SYNTHESIZED_WIRE_24);


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_37);



SYNTHESIZED_WIRE_1 <= NOT(SYNTHESIZED_WIRE_38);



SYNTHESIZED_WIRE_3 <= NOT(SYNTHESIZED_WIRE_36);



C <= SYNTHESIZED_WIRE_24 XOR SR;


V <= SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_27 XOR SR;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_28 XOR SR;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_29 XOR SR;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_38 XOR SR;


Z <= NOT(SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_36);


END bdf_type;