library verilog;
use verilog.vl_types.all;
entity ParteA_vlg_vec_tst is
end ParteA_vlg_vec_tst;
